bind wrap_fifo_c generic_twoport bind_fifo_c(.*);

